// megafunction wizard: %ALTLVDS%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altlvds_rx 

// ============================================================
// File Name: linki.v
// Megafunction Name(s):
// 			altlvds_rx
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.1 Build 350 03/24/2010 SP 2 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2010 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module linki (
	rx_in,
	rx_inclock,
	rx_reset,
	rx_dpa_locked,
	rx_locked,
	rx_out,
	rx_outclock);

	input	[8:0]  rx_in;
	input	  rx_inclock;
	input	[8:0]  rx_reset;
	output	[8:0]  rx_dpa_locked;
	output	  rx_locked;
	output	[35:0]  rx_out;
	output	  rx_outclock;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri0	[8:0]  rx_reset;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  sub_wire0;
	wire [35:0] sub_wire1;
	wire  sub_wire2;
	wire [8:0] sub_wire3;
	wire  rx_locked = sub_wire0;
	wire [35:0] rx_out = sub_wire1[35:0];
	wire  rx_outclock = sub_wire2;
	wire [8:0] rx_dpa_locked = sub_wire3[8:0];

	altlvds_rx	altlvds_rx_component (
				.rx_inclock (rx_inclock),
				.rx_reset (rx_reset),
				.rx_in (rx_in),
				.rx_locked (sub_wire0),
				.rx_out (sub_wire1),
				.rx_outclock (sub_wire2),
				.rx_dpa_locked (sub_wire3),
				.dpa_pll_cal_busy (),
				.dpa_pll_recal (1'b0),
				.pll_areset (1'b0),
				.pll_phasecounterselect (),
				.pll_phasedone (1'b1),
				.pll_phasestep (),
				.pll_phaseupdown (),
				.pll_scanclk (),
				.rx_cda_max (),
				.rx_cda_reset ({9{1'b0}}),
				.rx_channel_data_align ({9{1'b0}}),
				.rx_coreclk ({9{1'b1}}),
				.rx_data_align (1'b0),
				.rx_data_align_reset (1'b0),
				.rx_data_reset (1'b0),
				.rx_deskew (1'b0),
				.rx_divfwdclk (),
				.rx_dpa_lock_reset ({9{1'b0}}),
				.rx_dpll_enable ({9{1'b1}}),
				.rx_dpll_hold ({9{1'b0}}),
				.rx_dpll_reset ({9{1'b0}}),
				.rx_enable (1'b1),
				.rx_fifo_reset ({9{1'b0}}),
				.rx_pll_enable (1'b1),
				.rx_readclock (1'b0),
				.rx_syncclock (1'b0));
	defparam
		altlvds_rx_component.common_rx_tx_pll = "OFF",
		altlvds_rx_component.deserialization_factor = 4,
		altlvds_rx_component.enable_dpa_mode = "ON",
		altlvds_rx_component.implement_in_les = "OFF",
		altlvds_rx_component.inclock_period = 7813,
		altlvds_rx_component.input_data_rate = 512,
		altlvds_rx_component.intended_device_family = "Arria II GX",
		altlvds_rx_component.lpm_hint = "CBX_MODULE_PREFIX=linki",
		altlvds_rx_component.lpm_type = "altlvds_rx",
		altlvds_rx_component.number_of_channels = 9,
		altlvds_rx_component.outclock_resource = "AUTO",
		altlvds_rx_component.registered_output = "ON",
		altlvds_rx_component.use_external_pll = "OFF",
		altlvds_rx_component.enable_dpa_align_to_rising_edge_only = "OFF",
		altlvds_rx_component.enable_dpa_initial_phase_selection = "OFF";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: Bitslip NUMERIC "4"
// Retrieval info: PRIVATE: Channel_Data_Align_Max NUMERIC "0"
// Retrieval info: PRIVATE: Channel_Data_Align_Reset NUMERIC "0"
// Retrieval info: PRIVATE: Clock_Mode NUMERIC "0"
// Retrieval info: PRIVATE: Data_rate STRING "512"
// Retrieval info: PRIVATE: Deser_Factor NUMERIC "4"
// Retrieval info: PRIVATE: Dpa_Locked NUMERIC "1"
// Retrieval info: PRIVATE: Dpll_Enable NUMERIC "0"
// Retrieval info: PRIVATE: Dpll_Hold NUMERIC "0"
// Retrieval info: PRIVATE: Dpll_Reset NUMERIC "1"
// Retrieval info: PRIVATE: Enable_DPA_Mode STRING "ON"
// Retrieval info: PRIVATE: Ext_PLL STRING "OFF"
// Retrieval info: PRIVATE: Fifo_Reset NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
// Retrieval info: PRIVATE: Int_Device STRING "Arria II GX"
// Retrieval info: PRIVATE: LVDS_Mode NUMERIC "1"
// Retrieval info: PRIVATE: Le_Serdes STRING "OFF"
// Retrieval info: PRIVATE: Num_Channel NUMERIC "9"
// Retrieval info: PRIVATE: PLL_Enable NUMERIC "0"
// Retrieval info: PRIVATE: PLL_Freq STRING "128.00"
// Retrieval info: PRIVATE: PLL_Period STRING "7.813"
// Retrieval info: PRIVATE: Reg_InOut NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: Use_Clock_Resc STRING "AUTO"
// Retrieval info: PRIVATE: Use_Common_Rx_Tx_Plls NUMERIC "0"
// Retrieval info: PRIVATE: Use_Data_Align NUMERIC "0"
// Retrieval info: PRIVATE: Use_Lock NUMERIC "1"
// Retrieval info: PRIVATE: Use_Pll_Areset NUMERIC "0"
// Retrieval info: CONSTANT: COMMON_RX_TX_PLL STRING "OFF"
// Retrieval info: CONSTANT: DESERIALIZATION_FACTOR NUMERIC "4"
// Retrieval info: CONSTANT: ENABLE_DPA_MODE STRING "ON"
// Retrieval info: CONSTANT: IMPLEMENT_IN_LES STRING "OFF"
// Retrieval info: CONSTANT: INCLOCK_PERIOD NUMERIC "7813"
// Retrieval info: CONSTANT: INPUT_DATA_RATE NUMERIC "512"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altlvds_rx"
// Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "9"
// Retrieval info: CONSTANT: OUTCLOCK_RESOURCE STRING "AUTO"
// Retrieval info: CONSTANT: REGISTERED_OUTPUT STRING "ON"
// Retrieval info: CONSTANT: USE_EXTERNAL_PLL STRING "OFF"
// Retrieval info: CONSTANT: enable_dpa_align_to_rising_edge_only STRING "OFF"
// Retrieval info: CONSTANT: enable_dpa_initial_phase_selection STRING "OFF"
// Retrieval info: USED_PORT: rx_dpa_locked 0 0 9 0 OUTPUT NODEFVAL rx_dpa_locked[8..0]
// Retrieval info: USED_PORT: rx_in 0 0 9 0 INPUT NODEFVAL rx_in[8..0]
// Retrieval info: USED_PORT: rx_inclock 0 0 0 0 INPUT_CLK_EXT GND rx_inclock
// Retrieval info: USED_PORT: rx_locked 0 0 0 0 OUTPUT VCC rx_locked
// Retrieval info: USED_PORT: rx_out 0 0 36 0 OUTPUT NODEFVAL rx_out[35..0]
// Retrieval info: USED_PORT: rx_outclock 0 0 0 0 OUTPUT NODEFVAL rx_outclock
// Retrieval info: USED_PORT: rx_reset 0 0 9 0 INPUT GND rx_reset[8..0]
// Retrieval info: CONNECT: @rx_in 0 0 9 0 rx_in 0 0 9 0
// Retrieval info: CONNECT: rx_out 0 0 36 0 @rx_out 0 0 36 0
// Retrieval info: CONNECT: @rx_inclock 0 0 0 0 rx_inclock 0 0 0 0
// Retrieval info: CONNECT: rx_locked 0 0 0 0 @rx_locked 0 0 0 0
// Retrieval info: CONNECT: @rx_reset 0 0 9 0 rx_reset 0 0 9 0
// Retrieval info: CONNECT: rx_dpa_locked 0 0 9 0 @rx_dpa_locked 0 0 9 0
// Retrieval info: CONNECT: rx_outclock 0 0 0 0 @rx_outclock 0 0 0 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL linki.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL linki.ppf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL linki.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL linki.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL linki.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL linki_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL linki_bb.v FALSE
// Retrieval info: LIB_FILE: altera_mf
// Retrieval info: CBX_MODULE_PREFIX: ON
